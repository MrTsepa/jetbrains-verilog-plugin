module Foo (
	input foo
	);

endmodule
