module Biz (
	input biz
	);

endmodule
